mem[00]=32'h02000060;
mem[01]=32'h00807C2E;
mem[02]=32'hBC2E0001;
mem[03]=32'h00020000;
mem[04]=32'h00003C2F;
mem[05]=32'hFC2E0003;
mem[06]=32'h00040000;
mem[07]=32'h0000BC2E;
mem[08]=32'h00610005;
mem[09]=32'h00610A00;
mem[10]=32'h0060A400;
mem[11]=32'h7C20D200;
mem[12]=32'h020001FF;
mem[13]=32'h0100BC10;
mem[14]=32'h01FF7C20;
mem[15]=32'hBC100300;
mem[16]=32'h7C200100;
mem[17]=32'h020002FF;
mem[18]=32'h0100BC10;
mem[19]=32'h02FF7C20;
mem[20]=32'hBC100300;
mem[21]=32'h754E0100;
mem[22]=32'h01FF7C20;
mem[23]=32'h10100100;
mem[24]=32'h01000002;
mem[25]=32'h0061754E;
mem[26]=32'h0067F0FF;
mem[27]=32'h7C20FAFF;
mem[28]=32'h0001FFFF;
mem[29]=32'h754E1012;
mem[30]=32'h01FF7C20;
mem[31]=32'h10100100;
mem[32]=32'h02000002;
mem[33]=32'hF8FF0066;
mem[34]=32'h01FF7C20;
mem[35]=32'h81100000;
mem[36]=32'h7C20754E;
mem[37]=32'h010002FF;
mem[38]=32'h00021010;
mem[39]=32'h754E0100;
mem[40]=32'hF0FF0061;
mem[41]=32'hFAFF0067;
mem[42]=32'h02FF7C20;
mem[43]=32'h10120000;
mem[44]=32'h7C20754E;
mem[45]=32'h010002FF;
mem[46]=32'h00021010;
mem[47]=32'h00670200;
mem[48]=32'h7C20F8FF;
mem[49]=32'h000002FF;
mem[50]=32'h754E8110;
mem[51]=32'h4B003C12;
mem[52]=32'hA6FF0061;
mem[53]=32'hDCFF0061;
mem[54]=32'h36003C12;
mem[55]=32'h9AFF0061;
mem[56]=32'hD0FF0061;
mem[57]=32'h68003C12;
mem[58]=32'h8EFF0061;
mem[59]=32'hC4FF0061;
mem[60]=32'h0D003C12;
mem[61]=32'h82FF0061;
mem[62]=32'hB8FF0061;
mem[63]=32'h0061754E;
mem[64]=32'h006758FF;
mem[65]=32'h00610E00;
mem[66]=32'h00678AFF;
mem[67]=32'h00601400;
mem[68]=32'h0061EEFF;
mem[69]=32'h006152FF;
mem[70]=32'h00611800;
mem[71]=32'h754E96FF;
mem[72]=32'h7EFF0061;
mem[73]=32'h08000061;
mem[74]=32'h4EFF0061;
mem[75]=32'h754E754E;
mem[76]=32'h0000754E;
